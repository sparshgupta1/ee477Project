
* LOT: T26X                  WAF: 1011
* Temperature_parameters=Default
.MODEL TSMC20N NMOS (                                LEVEL   = 49
+VERSION = 3.1            TNOM    = 27             TOX     = 4.1E-9
+XJ      = 1E-7           NCH     = 2.3549E17      VTH0    = 0.3796589
+K1      = 0.5935169      K2      = 2.38533E-3     K3      = 1E-3
+K3B     = 3.1905105      W0      = 1E-7           NLX     = 1.786849E-7
+DVT0W   = 0              DVT1W   = 0              DVT2W   = 0
+DVT0    = 1.7203781      DVT1    = 0.4308344      DVT2    = 0.0467521
+U0      = 269.0634518    UA      = -1.188565E-9   UB      = 1.930877E-18
+UC      = 2.224818E-11   VSAT    = 9.67502E4      A0      = 2
+AGS     = 0.4169677      B0      = -1.063955E-8   B1      = -1E-7
+KETA    = -7.704208E-3   A1      = 7.99632E-4     A2      = 0.999873
+RDSW    = 105            PRWG    = 0.5            PRWB    = -0.2
+WR      = 1              WINT    = 2.025957E-9    LINT    = 1.028309E-8
+XL      = -2E-8          XW      = -1E-8          DWG     = -6.4982E-10
+DWB     = 1.217904E-8    VOFF    = -0.0901723     NFACTOR = 2.3820479
+CIT     = 0              CDSC    = 2.4E-4         CDSCD   = 0
+CDSCB   = 0              ETA0    = 1.448044E-3    ETAB    = -2.754731E-4
+DSUB    = 0.0110906      PCLM    = 1.0622551      PDIBLC1 = 0.3172281
+PDIBLC2 = 3.755701E-3    PDIBLCB = -0.1           DROUT   = 0.783102
+PSCBE1  = 5.995957E10    PSCBE2  = 5.686023E-8    PVAG    = 0.3568363
+DELTA   = 0.01           RSH     = 6.7            MOBMOD  = 1
+PRT     = 0              UTE     = -1.5           KT1     = -0.11
+KT1L    = 0              KT2     = 0.022          UA1     = 4.31E-9
+UB1     = -7.61E-18      UC1     = -5.6E-11       AT      = 3.3E4
+WL      = 0              WLN     = 1              WW      = 0
+WWN     = 1              WWL     = 0              LL      = 0
+LLN     = 1              LW      = 0              LWN     = 1
+LWL     = 0              CAPMOD  = 2              XPART   = 0.5
+CGDO    = 7.45E-10       CGSO    = 7.45E-10       CGBO    = 1E-12
+CJ      = 9.725136E-4    PB      = 0.7292509      MJ      = 0.3610145
+CJSW    = 2.269386E-10   PBSW    = 0.6351005      MJSW    = 0.1
+CJSWG   = 3.3E-10        PBSWG   = 0.6351005      MJSWG   = 0.1
+CF      = 0              PVTH0   = -2.139932E-3   PRDSW   = -1.2311975
+PK2     = 1.860342E-3    WKETA   = 1.76355E-3     LKETA   = -5.667186E-3
+PU0     = -0.2295277     PUA     = -2.87112E-11   PUB     = 0
+PVSAT   = 1.427606E3     PETA0   = 1E-4           PKETA   = -1.196986E-3    )



* LOT: T26X                  WAF: 1011
* Temperature_parameters=Default
.MODEL TSMC20P PMOS (                                LEVEL   = 49
+VERSION = 3.1            TNOM    = 27             TOX     = 4.1E-9
+XJ      = 1E-7           NCH     = 4.1589E17      VTH0    = -0.4215645
+K1      = 0.5955538      K2      = 0.0265154      K3      = 0
+K3B     = 10.7990376     W0      = 1E-6           NLX     = 7.393151E-8
+DVT0W   = 0              DVT1W   = 0              DVT2W   = 0
+DVT0    = 0.3622323      DVT1    = 0.2560341      DVT2    = 0.1
+U0      = 119.2085214    UA      = 1.656038E-9    UB      = 1E-21
+UC      = -1E-10         VSAT    = 1.840486E5     A0      = 1.7659056
+AGS     = 0.4199318      B0      = 9.960505E-7    B1      = 3.37199E-6
+KETA    = 0.0126497      A1      = 0.4537105      A2      = 0.3
+RDSW    = 201.0196067    PRWG    = 0.5            PRWB    = -0.5
+WR      = 1              WINT    = 0              LINT    = 2.42201E-8
+XL      = -2E-8          XW      = -1E-8          DWG     = -2.790988E-8
+DWB     = 5.977646E-9    VOFF    = -0.1035186     NFACTOR = 1.8044589
+CIT     = 0              CDSC    = 2.4E-4         CDSCD   = 0
+CDSCB   = 0              ETA0    = 0.0079869      ETAB    = -0.115204
+DSUB    = 0.940025       PCLM    = 1.9711817      PDIBLC1 = 0
+PDIBLC2 = 0.0195957      PDIBLCB = -1E-3          DROUT   = 5.830459E-4
+PSCBE1  = 2.224265E9     PSCBE2  = 6.4242E-10     PVAG    = 10.2269693
+DELTA   = 0.01           RSH     = 7.6            MOBMOD  = 1
+PRT     = 0              UTE     = -1.5           KT1     = -0.11
+KT1L    = 0              KT2     = 0.022          UA1     = 4.31E-9
+UB1     = -7.61E-18      UC1     = -5.6E-11       AT      = 3.3E4
+WL      = 0              WLN     = 1              WW      = 0
+WWN     = 1              WWL     = 0              LL      = 0
+LLN     = 1              LW      = 0              LWN     = 1
+LWL     = 0              CAPMOD  = 2              XPART   = 0.5
+CGDO    = 6.52E-10       CGSO    = 6.52E-10       CGBO    = 1E-12
+CJ      = 1.156829E-3    PB      = 0.8604313      MJ      = 0.4161985
+CJSW    = 1.800318E-10   PBSW    = 0.6161205      MJSW    = 0.2735145
+CJSWG   = 4.22E-10       PBSWG   = 0.6161205      MJSWG   = 0.2735145
+CF      = 0              PVTH0   = 1.121114E-3    PRDSW   = 12.2644118
+PK2     = 1.671328E-3    WKETA   = 2.478808E-3    LKETA   = -2.85111E-3
+PU0     = -1.8187729     PUA     = -7.23748E-11   PUB     = 1E-21
+PVSAT   = -50            PETA0   = 1E-4           PKETA   = 2.650105E-3     )

